** Profile: "SCHEMATIC1-iranpour-p1"  [ C:\Users\ZahraIranpour\Desktop\term 6\elec sanati\hw\shabih sazi\project1-SCHEMATIC1-iranpour-p1.sim ] 

** Creating circuit file "project1-SCHEMATIC1-iranpour-p1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 75ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\project1-SCHEMATIC1.net" 


.END
